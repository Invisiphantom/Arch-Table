`ifndef CONFIG_SV
`define CONFIG_SV

package config_pkg;
	// parameters
	parameter AXI_BURST_NUM = 16;


	
endpackage

`endif
